module sys

#flag darwin -framework OpenGL
